library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity cpu is
end cpu;

architecture Behavioral of cpu is
	component pop_cpu
		port ( outRam2OE : out STD_LOGIC; 
    RAM1WE : out STD_LOGIC; 
    outRam2WE : out STD_LOGIC; 
    outwdn : out STD_LOGIC; 
    outrdn : out STD_LOGIC; 
    RAM1EN : out STD_LOGIC; 
    tsre : in STD_LOGIC := 'X'; 
    outRam2EN : out STD_LOGIC; 
    RAM1OE : out STD_LOGIC; 
    dataReady : in STD_LOGIC := 'X'; 
    inclk : in STD_LOGIC := 'X'; 
    RAM1data : inout STD_LOGIC_VECTOR ( 15 downto 0 ); 
    outRam2Data : inout STD_LOGIC_VECTOR ( 15 downto 0 ); 
    l7 : out STD_LOGIC_VECTOR ( 6 downto 0 ); 
    r7 : out STD_LOGIC_VECTOR ( 6 downto 0 ); 
    RAM1addr : out STD_LOGIC_VECTOR ( 17 downto 0 ); 
    ins : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    outRam2Addr : out STD_LOGIC_VECTOR ( 17 downto 0 ));
	end component;
	signal clk : std_logic := '1';
	signal RAM1OE : STD_LOGIC := '0';
	signal RAM1WE : STD_LOGIC := '0';
	signal RAM1EN : STD_LOGIC := '0';
	signal RAM1addr : STD_LOGIC_VECTOR (17 downto 0) :=(others=>'0');
	signal RAM1data : STD_LOGIC_VECTOR (15 downto 0) :=(others=>'0');
	signal Ram2OE : STD_LOGIC := '0';
	signal Ram2WE : STD_LOGIC := '0';
	signal Ram2EN : STD_LOGIC := '0';
	signal Ram2Addr : STD_LOGIC_VECTOR(17 downto 0) :=(others=>'0');
	signal Ram2Data : STD_LOGIC_VECTOR(15 downto 0) :=(others=>'0');
	signal dataReady : STD_LOGIC := '0';
	signal tsre : STD_LOGIC := '0';
	signal rdn : STD_LOGIC := '0';
	signal wdn : STD_LOGIC := '0';
	signal cnt : STD_LOGIC_VECTOR(3 downto 0) := "0000";
begin
	c : pop_cpu port map(inclk => clk, RAM1OE => RAM1OE, RAM1WE => RAM1WE, RAM1EN => RAM1EN, RAM1addr => RAM1addr, RAM1data => RAM1Data,
				outRam2OE => Ram2OE, outRam2WE => RAM2WE, outRam2EN => RAM2EN, outRam2Addr => Ram2Addr, outRam2Data => RAM2Data,
				dataReady => dataready, tsre =>tsre, outrdn=>rdn, outwdn=>wdn);
	clk <= not clk after 100ns;
	cnt <= cnt + "1" after 200ns;
	process(Ram2Addr, RAM2Data)
	begin
	case Ram2Addr is
		when "00"&X"0000" =>
			Ram2Data <= X"0000" after 10ns;
		when "00"&X"0001" =>
			Ram2Data <= X"0000"  after 10ns;
		when "00"&X"0002" =>
			Ram2Data <= X"0800" after 10ns;
		when "00"&X"0003" =>
			Ram2Data <= X"1044" after 10ns;


		when "00"&X"0048" =>
			Ram2Data <= X"6807" after 10ns;
		when "00"&X"0049" =>
			Ram2Data <= X"F001" after 10ns;
		when "00"&X"004A" =>
			Ram2Data <= X"68BF" after 10ns;
		when "00"&X"004B" =>
			Ram2Data <= X"3000" after 10ns;
		when "00"&X"004C" =>
			Ram2Data <= X"4810" after 10ns;
		when "00"&X"004D" =>
			Ram2Data <= X"6400" after 10ns;
		when "00"&X"004E" =>
			Ram2Data <= X"0800" after 10ns;
		when "00"&X"004F" =>
			Ram2Data <= X"6EBF" after 10ns;
		when "00"&X"0050" =>
			Ram2Data <= X"36C0" after 10ns;
		when "00"&X"0051" =>
			Ram2Data <= X"4E10" after 10ns;
		when "00"&X"0052" =>
			Ram2Data <= X"6800" after 10ns;
		when "00"&X"0053" =>
			Ram2Data <= X"DE00" after 10ns;
		when "00"&X"0054" =>
			Ram2Data <= X"DE01" after 10ns;
		when "00"&X"0055" =>
			Ram2Data <= X"DE02" after 10ns;
		when "00"&X"0056" =>
			Ram2Data <= X"DE03" after 10ns;
		when "00"&X"0057" =>
			Ram2Data <= X"DE04" after 10ns;
		when "00"&X"0058" =>
			Ram2Data <= X"DE05" after 10ns;
		when "00"&X"0059" =>
			Ram2Data <= X"EF40" after 10ns;
		when "00"&X"005A" =>
			Ram2Data <= X"4F03" after 10ns;
		when "00"&X"005B" =>
			Ram2Data <= X"0800" after 10ns;
		when "00"&X"005C" =>
			Ram2Data <= X"104A" after 10ns;
		when "00"&X"005D" =>
			Ram2Data <= X"6EBF" after 10ns;
		when "00"&X"005E" =>
			Ram2Data <= X"36C0" after 10ns;
		when "00"&X"005F" =>
			Ram2Data <= X"684F" after 10ns;
		when "00"&X"0060" =>
			Ram2Data <= X"DE00" after 10ns;
		when "00"&X"0061" =>
			Ram2Data <= X"0800" after 10ns;
		when "00"&X"0062" =>
			Ram2Data <= X"EF40" after 10ns;


		when "00"&X"00A7" =>
			Ram2Data <= X"0800";
		when "00"&X"00A8" =>
			Ram2Data <= X"6EBF";
		when "00"&X"00A9" =>
			Ram2Data <= X"36C0";
		when "00"&X"00AA" =>
			Ram2Data <= X"4E01";
		when "00"&X"00AB" =>
			Ram2Data <= X"9E00";
		when "00"&X"00AC" =>
			Ram2Data <= X"6E01";
		when "00"&X"00AD" =>
			Ram2Data <= X"E8CC";
		when "00"&X"00AE" =>
			Ram2Data <= X"20F8";
		when "00"&X"00AF" =>
			Ram2Data <= X"0800";
		when "00"&X"00B0" =>
			Ram2Data <= X"EF00";
		when "00"&X"00B1" =>
			Ram2Data <= X"0800";

		--when "000000000000000100" =>
			--Ram2Data <= "0110100000100000"; 
		--when "000000000000000101" =>
			--Ram2Data <= X"db20";
		--when "000000000000000110" =>
			--Ram2Data <= X"db41"; 
		--when "000000000000000111" =>
			--Ram2Data <= X"e145";

		--when "000000000000001000" =>
			--Ram2Data <= X"e149";	 
		--when "000000000000001001" =>
			--Ram2Data <= X"4b02";
		--when "000000000000001010" =>
			--Ram2Data <= X"4cff";
		--when "000000000000001011" =>
			--Ram2Data <= X"2cf9"; 

		when others => 
			Ram2Data <= "0000100000000000"; --nop
	end case;
	end process;
	process(RAM1addr,rdn)
	begin
		if(RAM1EN='0' and RAM1WE='1')then
			case RAM1addr is
				when "00"&X"BF00" =>
					RAM1data <= X"1001";
				when others =>
					RAM1data <= X"0000";
			end case;
		else
			if(rdn='0')then
				RAM1data <= X"1001";
			end if;
			dataReady <= '1';
			tsre <= '1';
		end if;
	end process;
end Behavioral;